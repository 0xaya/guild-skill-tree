No,スキル名,系統,タイプ,説明,必要ランク,ギルドコイン,記憶の書,剛力Ⅰ,剛力Ⅱ,剛力Ⅲ,鉄壁Ⅰ,鉄壁Ⅱ,鉄壁Ⅲ,魔道Ⅰ,魔道Ⅱ,魔道Ⅲ,精微Ⅰ,精微Ⅱ,精微Ⅲ,疾風Ⅰ,疾風Ⅱ,疾風Ⅲ,救済Ⅰ,救済Ⅱ,救済Ⅲ
11,腕力ⅠLv1,腕力系統,パッシブ,腕力を1%増加,2,10,,,,,,,,,,,,,,,,,,,
11,腕力ⅠLv2,腕力系統,パッシブ,腕力を2%増加,3,30,,,,,,,,,,,,,,,,,,,
11,腕力ⅠLv3,腕力系統,パッシブ,腕力を4%増加,4,80,10,20,,,,,,,,,,,,,,,,,
11,腕力ⅠLv4,腕力系統,パッシブ,腕力を7%増加,5,140,20,20,10,,,,,,,,,,,,,,,,
11,腕力ⅠLv5,腕力系統,パッシブ,腕力を10%増加,6,250,30,20,20,10,,,,,,,,,,,,,,,
12,体力ⅠLv1,体力系統,パッシブ,体力を1%増加,2,10,,,,,,,,,,,,,,,,,,,
12,体力ⅠLv2,体力系統,パッシブ,体力を2%増加,3,30,,,,,,,,,,,,,,,,,,,
12,体力ⅠLv3,体力系統,パッシブ,体力を4%増加,4,80,10,,,,20,,,,,,,,,,,,,,
12,体力ⅠLv4,体力系統,パッシブ,体力を7%増加,5,140,20,,,,20,10,,,,,,,,,,,,,
12,体力ⅠLv5,体力系統,パッシブ,体力を10%増加,6,250,30,,,,20,20,10,,,,,,,,,,,,
13,速さⅠLv1,速さ系統,パッシブ,速さを1%増加,2,10,,,,,,,,,,,,,,,,,,,
13,速さⅠLv2,速さ系統,パッシブ,速さを2%増加,3,30,,,,,,,,,,,,,,,,,,,
13,速さⅠLv3,速さ系統,パッシブ,速さを4%増加,4,80,10,,,,,,,,,,,,,20,,,,,
13,速さⅠLv4,速さ系統,パッシブ,速さを7%増加,5,140,20,,,,,,,,,,,,,20,10,,,,
13,速さⅠLv5,速さ系統,パッシブ,速さを10%増加,6,250,30,,,,,,,,,,,,,20,20,10,,,
14,知力ⅠLv1,知力系統,パッシブ,知力を1%増加,2,10,,,,,,,,,,,,,,,,,,,
14,知力ⅠLv2,知力系統,パッシブ,知力を2%増加,3,30,,,,,,,,,,,,,,,,,,,
14,知力ⅠLv3,知力系統,パッシブ,知力を4%増加,4,80,10,,,,,,,20,,,,,,,,,,,
14,知力ⅠLv4,知力系統,パッシブ,知力を7%増加,5,140,20,,,,,,,20,10,,,,,,,,,,
14,知力ⅠLv5,知力系統,パッシブ,知力を10%増加,6,250,30,,,,,,,20,20,10,,,,,,,,,
15,器用ⅠLv1,器用系統,パッシブ,器用を1%増加,2,10,,,,,,,,,,,,,,,,,,,
15,器用ⅠLv2,器用系統,パッシブ,器用を2%増加,3,30,,,,,,,,,,,,,,,,,,,
15,器用ⅠLv3,器用系統,パッシブ,器用を4%増加,4,80,10,,,,,,,,,,20,,,,,,,,
15,器用ⅠLv4,器用系統,パッシブ,器用を7%増加,5,140,20,,,,,,,,,,20,10,,,,,,,
15,器用ⅠLv5,器用系統,パッシブ,器用を10%増加,6,250,30,,,,,,,,,,20,20,10,,,,,,
16,精神ⅠLv1,精神系統,パッシブ,精神を1%増加,2,10,,,,,,,,,,,,,,,,,,,
16,精神ⅠLv2,精神系統,パッシブ,精神を2%増加,3,30,,,,,,,,,,,,,,,,,,,
16,精神ⅠLv3,精神系統,パッシブ,精神を4%増加,4,80,10,,,,,,,,,,,,,,,,20,,
16,精神ⅠLv4,精神系統,パッシブ,精神を7%増加,5,140,20,,,,,,,,,,,,,,,,20,10,
16,精神ⅠLv5,精神系統,パッシブ,精神を10%増加,6,250,30,,,,,,,,,,,,,,,,20,20,10
21,HPⅡLv1,腕力系統,パッシブ,最大HPを2%増加,3,12,,,,,,,,,,,,,,,,,,,
21,HPⅡLv2,腕力系統,パッシブ,最大HPを4%増加,4,36,10,20,,,,,,,,,,,,,,,,,
21,HPⅡLv3,腕力系統,パッシブ,最大HPを6%増加,5,96,20,40,,,,,,,,,,,,,,,,,
21,HPⅡLv4,腕力系統,パッシブ,最大HPを9%増加,6,168,40,40,20,,,,,,,,,,,,,,,,
21,HPⅡLv5,腕力系統,パッシブ,最大HPを12%増加,7,300,60,40,20,20,,,,,,,,,,,,,,,
212,物理クリティカル発動率ⅡLv1,腕力系統,パッシブ,物理クリティカル発動率を1%増加,4,12,,,,,,,,,,,,,,,,,,,
212,物理クリティカル発動率ⅡLv2,腕力系統,パッシブ,物理クリティカル発動率を2%増加,5,36,10,20,,,,,,,,,,,,,,,,,
212,物理クリティカル発動率ⅡLv3,腕力系統,パッシブ,物理クリティカル発動率を4%増加,6,96,20,40,,,,,,,,,,,,,,,,,
212,物理クリティカル発動率ⅡLv4,腕力系統,パッシブ,物理クリティカル発動率を7%増加,7,168,40,40,20,,,,,,,,,,,,,,,,
212,物理クリティカル発動率ⅡLv5,腕力系統,パッシブ,物理クリティカル発動率を10%増加,8,300,60,40,20,20,,,,,,,,,,,,,,,
31,攻撃速度ⅢLv1,腕力系統,パッシブ,攻撃速度を5%増加,6,30,,,,,,,,,,,,,,,,,,,
31,攻撃速度ⅢLv2,腕力系統,パッシブ,攻撃速度を10%増加,7,80,20,40,,,,,,,,,,,,,,,,,
31,攻撃速度ⅢLv3,腕力系統,パッシブ,攻撃速度を15%増加,8,140,40,40,20,,,,,,,,,,,,,,,,
31,攻撃速度ⅢLv4,腕力系統,パッシブ,攻撃速度を20%増加,9,250,80,40,20,20,,,,,,,,,,,,,,,
31,攻撃速度ⅢLv5,腕力系統,パッシブ,攻撃速度を30%増加,10,400,120,80,40,20,,,,,,,,,,,,,,,
323,腕力ⅡLv1,腕力系統,パッシブ,腕力を2%増加,7,30,,,,,,,,,,,,,,,,,,,
323,腕力ⅡLv2,腕力系統,パッシブ,腕力を4%増加,8,80,20,40,,,,,,,,,,,,,,,,,
323,腕力ⅡLv3,腕力系統,パッシブ,腕力を6%増加,9,140,40,40,20,,,,,,,,,,,,,,,,
323,腕力ⅡLv4,腕力系統,パッシブ,腕力を10%増加,10,250,80,40,20,20,,,,,,,,,,,,,,,
323,腕力ⅡLv5,腕力系統,パッシブ,腕力を15%増加,11,400,120,80,40,20,,,,,,,,,,,,,,,
324,物理スキル威力ⅡLv1,腕力系統,パッシブ,物理スキル威力を1.05倍する,8,30,,,,,,,,,,,,,,,,,,,
324,物理スキル威力ⅡLv2,腕力系統,パッシブ,物理スキル威力を1.10倍する,9,80,20,40,,,,,,,,,,,,,,,,,
324,物理スキル威力ⅡLv3,腕力系統,パッシブ,物理スキル威力を1.15倍する,10,140,40,40,20,,,,,,,,,,,,,,,,
324,物理スキル威力ⅡLv4,腕力系統,パッシブ,物理スキル威力を1.20倍する,11,250,80,40,20,20,,,,,,,,,,,,,,,
324,物理スキル威力ⅡLv5,腕力系統,パッシブ,物理スキル威力を1.25倍する,12,400,120,80,40,20,,,,,,,,,,,,,,,
322,無双Lv1,腕力系統,アクティブ,詠唱時間1.5倍に増えて物理スキル威力1.2倍,10,50,50,,,,,,,,,,,,,,,,,,
322,無双Lv2,腕力系統,アクティブ,詠唱時間1.5倍に増えて物理スキル威力1.4倍,11,100,100,50,,,,,,,,,,,,,,,,,
322,無双Lv3,腕力系統,アクティブ,詠唱時間1.35倍に増えて物理スキル威力1.6倍,12,180,150,60,30,,,,,,,,,,,,,,,,
322,無双Lv4,腕力系統,アクティブ,詠唱時間1.35倍に増えて物理スキル威力1.8倍,13,300,200,70,40,20,,,,,,,,,,,,,,,
322,無双Lv5,腕力系統,アクティブ,詠唱時間1.25倍に増えて物理スキル威力2.0倍,14,450,250,80,50,30,,,,,,,,,,,,,,,
23,防御力ⅠLv1,体力系統,パッシブ,防御力を2%増加,3,12,,,,,,,,,,,,,,,,,,,
23,防御力ⅠLv2,体力系統,パッシブ,防御力を4%増加,4,36,10,,,,20,,,,,,,,,,,,,,
23,防御力ⅠLv3,体力系統,パッシブ,防御力を6%増加,5,96,20,,,,40,,,,,,,,,,,,,,
23,防御力ⅠLv4,体力系統,パッシブ,防御力を9%増加,6,168,40,,,,40,20,,,,,,,,,,,,,
23,防御力ⅠLv5,体力系統,パッシブ,防御力を12%増加,7,300,60,,,,40,20,20,,,,,,,,,,,,
22,HPⅠLv1,体力系統,パッシブ,最大HPを2%増加,4,12,,,,,,,,,,,,,,,,,,,
22,HPⅠLv2,体力系統,パッシブ,最大HPを4%増加,5,36,10,,,,20,,,,,,,,,,,,,,
22,HPⅠLv3,体力系統,パッシブ,最大HPを6%増加,6,96,20,,,,40,,,,,,,,,,,,,,
22,HPⅠLv4,体力系統,パッシブ,最大HPを9%増加,7,168,40,,,,40,20,,,,,,,,,,,,,
22,HPⅠLv5,体力系統,パッシブ,最大HPを12%増加,8,300,60,,,,40,20,20,,,,,,,,,,,,
35,MPⅡLv1,体力系統,パッシブ,最大MPを3%増加,6,30,,,,,,,,,,,,,,,,,,,
35,MPⅡLv2,体力系統,パッシブ,最大MPを6%増加,7,80,20,,,,40,,,,,,,,,,,,,,
35,MPⅡLv3,体力系統,パッシブ,最大MPを10%増加,8,140,40,,,,40,20,,,,,,,,,,,,,
35,MPⅡLv4,体力系統,パッシブ,最大MPを15%増加,9,250,80,,,,40,20,20,,,,,,,,,,,,
35,MPⅡLv5,体力系統,パッシブ,最大MPを20%増加,10,400,120,,,,80,40,20,,,,,,,,,,,,
32,体力ⅡLv1,体力系統,パッシブ,体力を2%増加,7,30,,,,,,,,,,,,,,,,,,,
32,体力ⅡLv2,体力系統,パッシブ,体力を4%増加,8,80,20,,,,40,,,,,,,,,,,,,,
32,体力ⅡLv3,体力系統,パッシブ,体力を6%増加,9,140,40,,,,40,20,,,,,,,,,,,,,
32,体力ⅡLv4,体力系統,パッシブ,体力を10%増加,10,250,80,,,,40,20,20,,,,,,,,,,,,
32,体力ⅡLv5,体力系統,パッシブ,体力を15%増加,11,400,120,,,,80,40,20,,,,,,,,,,,,
34,EXP獲得率Lv1,体力系統,パッシブ,EXP獲得率を1.1倍する,8,30,,,,,,,,,,,,,,,,,,,
34,EXP獲得率Lv2,体力系統,パッシブ,EXP獲得率を1.15倍する,9,80,20,,,,40,,,,,,,,,,,,,,
34,EXP獲得率Lv3,体力系統,パッシブ,EXP獲得率を1.20倍する,10,140,40,,,,40,20,,,,,,,,,,,,,
34,EXP獲得率Lv4,体力系統,パッシブ,EXP獲得率を1.25倍する,11,250,80,,,,40,20,20,,,,,,,,,,,,
34,EXP獲得率Lv5,体力系統,パッシブ,EXP獲得率を1.30倍する,12,400,120,,,,80,40,20,,,,,,,,,,,,
33,不死Lv1,体力系統,アクティブ,MP半分消費してリヴァイブ（蘇生時HP20%）,10,50,50,,,,,,,,,,,,,,,,,,
33,不死Lv2,体力系統,アクティブ,MP半分消費してリヴァイブ（蘇生時HP40%）,11,100,100,,,,50,,,,,,,,,,,,,,
33,不死Lv3,体力系統,アクティブ,MP半分消費してリヴァイブ（蘇生時HP60%）,12,180,150,,,,60,30,,,,,,,,,,,,,
33,不死Lv4,体力系統,アクティブ,MP半分消費してリヴァイブ（蘇生時HP80%）,13,300,200,,,,70,40,20,,,,,,,,,,,,
33,不死Lv5,体力系統,アクティブ,MP半分消費してリヴァイブ（蘇生時HP100%）,14,450,250,,,,80,50,30,,,,,,,,,,,,
25,攻撃速度ⅠLv1,速さ系統,パッシブ,攻撃速度を3%増加,3,12,,,,,,,,,,,,,,,,,,,
25,攻撃速度ⅠLv2,速さ系統,パッシブ,攻撃速度を6%増加,4,36,10,,,,,,,,,,,,,20,,,,,
25,攻撃速度ⅠLv3,速さ系統,パッシブ,攻撃速度を10%増加,5,96,20,,,,,,,,,,,,,40,,,,,
25,攻撃速度ⅠLv4,速さ系統,パッシブ,攻撃速度を15%増加,6,168,40,,,,,,,,,,,,,40,20,,,,
25,攻撃速度ⅠLv5,速さ系統,パッシブ,攻撃速度を20%増加,7,300,60,,,,,,,,,,,,,40,20,20,,,
24,物理スキル威力ⅠLv1,速さ系統,パッシブ,物理スキル威力を1.03倍する,4,12,,,,,,,,,,,,,,,,,,,
24,物理スキル威力ⅠLv2,速さ系統,パッシブ,物理スキル威力を1.06倍する,5,36,10,,,,,,,,,,,,,20,,,,,
24,物理スキル威力ⅠLv3,速さ系統,パッシブ,物理スキル威力を1.09倍する,6,96,20,,,,,,,,,,,,,40,,,,,
24,物理スキル威力ⅠLv4,速さ系統,パッシブ,物理スキル威力を1.12倍する,7,168,40,,,,,,,,,,,,,40,20,,,,
24,物理スキル威力ⅠLv5,速さ系統,パッシブ,物理スキル威力を1.15倍する,8,300,60,,,,,,,,,,,,,40,20,20,,,
39,防御力ⅡLv1,速さ系統,パッシブ,防御力を3%増加,6,30,,,,,,,,,,,,,,,,,,,
39,防御力ⅡLv2,速さ系統,パッシブ,防御力を6%増加,7,80,20,,,,,,,,,,,,,40,,,,,
39,防御力ⅡLv3,速さ系統,パッシブ,防御力を9%増加,8,140,40,,,,,,,,,,,,,40,20,,,,
39,防御力ⅡLv4,速さ系統,パッシブ,防御力を13%増加,9,250,80,,,,,,,,,,,,,40,20,20,,,
39,防御力ⅡLv5,速さ系統,パッシブ,防御力を18%増加,10,400,120,,,,,,,,,,,,,80,40,20,,,
36,速さⅡLv1,速さ系統,パッシブ,速さを2%増加,7,30,,,,,,,,,,,,,,,,,,,
36,速さⅡLv2,速さ系統,パッシブ,速さを4%増加,8,80,20,,,,,,,,,,,,,40,,,,,
36,速さⅡLv3,速さ系統,パッシブ,速さを6%増加,9,140,40,,,,,,,,,,,,,40,20,,,,
36,速さⅡLv4,速さ系統,パッシブ,速さを10%増加,10,250,80,,,,,,,,,,,,,40,20,20,,,
36,速さⅡLv5,速さ系統,パッシブ,速さを15%増加,11,400,120,,,,,,,,,,,,,80,40,20,,,
38,詠唱速度ⅡLv1,速さ系統,パッシブ,詠唱速度を1.05倍する,8,30,,,,,,,,,,,,,,,,,,,
38,詠唱速度ⅡLv2,速さ系統,パッシブ,詠唱速度を1.10倍する,9,80,20,,,,,,,,,,,,,40,,,,,
38,詠唱速度ⅡLv3,速さ系統,パッシブ,詠唱速度を1.15倍する,10,140,40,,,,,,,,,,,,,40,20,,,,
38,詠唱速度ⅡLv4,速さ系統,パッシブ,詠唱速度を1.20倍する,11,250,80,,,,,,,,,,,,,40,20,20,,,
38,詠唱速度ⅡLv5,速さ系統,パッシブ,詠唱速度を1.25倍する,12,400,120,,,,,,,,,,,,,80,40,20,,,
37,明鏡Lv1,速さ系統,アクティブ,HP→MPに変換（HP10%消費してMP5%回復）,10,50,50,,,,,,,,,,,,,,,,,,
37,明鏡Lv2,速さ系統,アクティブ,HP→MPに変換（HP15%消費してMP10%回復）,11,100,100,,,,,,,,,,,,,50,,,,,
37,明鏡Lv3,速さ系統,アクティブ,HP→MPに変換（HP20%消費してMP15%回復）,12,180,150,,,,,,,,,,,,,60,30,,,,
37,明鏡Lv4,速さ系統,アクティブ,HP→MPに変換（HP25%消費してMP20%回復）,13,300,200,,,,,,,,,,,,,70,40,20,,,
37,明鏡Lv5,速さ系統,アクティブ,HP→MPに変換（HP30%消費してMP25%回復）,14,450,250,,,,,,,,,,,,,80,50,30,,,
27,魔法スキル威力ⅠLv1,知力系統,パッシブ,魔法スキル威力を1.05倍する,3,12,,,,,,,,,,,,,,,,,,,
27,魔法スキル威力ⅠLv2,知力系統,パッシブ,魔法スキル威力を1.10倍する,4,36,10,,,,,,,20,,,,,,,,,,,
27,魔法スキル威力ⅠLv3,知力系統,パッシブ,魔法スキル威力を1.15倍する,5,96,20,,,,,,,40,,,,,,,,,,,
27,魔法スキル威力ⅠLv4,知力系統,パッシブ,魔法スキル威力を1.20倍する,6,168,40,,,,,,,40,20,,,,,,,,,,
27,魔法スキル威力ⅠLv5,知力系統,パッシブ,魔法スキル威力を1.25倍する,7,300,60,,,,,,,40,20,20,,,,,,,,,
313,MPⅢLv1,知力系統,パッシブ,最大MPを3%増加,4,12,,,,,,,,,,,,,,,,,,,
313,MPⅢLv2,知力系統,パッシブ,最大MPを6%増加,5,36,10,,,,,,,20,,,,,,,,,,,
313,MPⅢLv3,知力系統,パッシブ,最大MPを10%増加,6,96,20,,,,,,,40,,,,,,,,,,,
313,MPⅢLv4,知力系統,パッシブ,最大MPを15%増加,7,168,40,,,,,,,40,20,,,,,,,,,,
313,MPⅢLv5,知力系統,パッシブ,最大MPを20%増加,8,300,60,,,,,,,40,20,20,,,,,,,,,
26,HPⅢLv1,知力系統,パッシブ,最大HPを2%増加,6,30,,,,,,,,,,,,,,,,,,,
26,HPⅢLv2,知力系統,パッシブ,最大HPを4%増加,7,80,20,,,,,,,40,,,,,,,,,,,
26,HPⅢLv3,知力系統,パッシブ,最大HPを6%増加,8,140,40,,,,,,,40,20,,,,,,,,,,
26,HPⅢLv4,知力系統,パッシブ,最大HPを9%増加,9,250,80,,,,,,,40,20,20,,,,,,,,,
26,HPⅢLv5,知力系統,パッシブ,最大HPを12%増加,10,400,120,,,,,,,80,40,20,,,,,,,,,
312,知力ⅡLv1,知力系統,パッシブ,知力を2%増加,7,30,,,,,,,,,,,,,,,,,,,
312,知力ⅡLv2,知力系統,パッシブ,知力を4%増加,8,80,20,,,,,,,40,,,,,,,,,,,
312,知力ⅡLv3,知力系統,パッシブ,知力を6%増加,9,140,40,,,,,,,40,20,,,,,,,,,,
312,知力ⅡLv4,知力系統,パッシブ,知力を10%増加,10,250,80,,,,,,,40,20,20,,,,,,,,,
312,知力ⅡLv5,知力系統,パッシブ,知力を15%増加,11,400,120,,,,,,,80,40,20,,,,,,,,,
310,魔法スキル威力ⅡLv1,知力系統,パッシブ,魔法スキル威力を1.08倍する,8,30,,,,,,,,,,,,,,,,,,,
310,魔法スキル威力ⅡLv2,知力系統,パッシブ,魔法スキル威力を1.16倍する,9,80,20,,,,,,,40,,,,,,,,,,,
310,魔法スキル威力ⅡLv3,知力系統,パッシブ,魔法スキル威力を1.24倍する,10,140,40,,,,,,,40,20,,,,,,,,,,
310,魔法スキル威力ⅡLv4,知力系統,パッシブ,魔法スキル威力を1.32倍する,11,250,80,,,,,,,40,20,20,,,,,,,,,
310,魔法スキル威力ⅡLv5,知力系統,パッシブ,魔法スキル威力を1.40倍する,12,400,120,,,,,,,80,40,20,,,,,,,,,
311,深淵Lv1,知力系統,アクティブ,1分間魔法スキルの威力を10%アップする,10,50,50,,,,,,,,,,,,,,,,,,
311,深淵Lv2,知力系統,アクティブ,1分間魔法スキルの威力を20%アップする,11,100,100,,,,,,,50,,,,,,,,,,,
311,深淵Lv3,知力系統,アクティブ,1分間魔法スキルの威力を30%アップする,12,180,150,,,,,,,60,30,,,,,,,,,,
311,深淵Lv4,知力系統,アクティブ,1分間魔法スキルの威力を40%アップする,13,300,200,,,,,,,70,40,20,,,,,,,,,
311,深淵Lv5,知力系統,アクティブ,1分間魔法スキルの威力を50%アップする,14,450,250,,,,,,,80,50,30,,,,,,,,,
29,物理クリティカル発動率ⅠLv1,器用系統,パッシブ,物理クリティカル発動率を1%増加,3,12,,,,,,,,,,,,,,,,,,,
29,物理クリティカル発動率ⅠLv2,器用系統,パッシブ,物理クリティカル発動率を2%増加,4,36,10,,,,,,,,,,20,,,,,,,,
29,物理クリティカル発動率ⅠLv3,器用系統,パッシブ,物理クリティカル発動率を4%増加,5,96,20,,,,,,,,,,40,,,,,,,,
29,物理クリティカル発動率ⅠLv4,器用系統,パッシブ,物理クリティカル発動率を7%増加,6,168,40,,,,,,,,,,40,20,,,,,,,
29,物理クリティカル発動率ⅠLv5,器用系統,パッシブ,物理クリティカル発動率を10%増加,7,300,60,,,,,,,,,,40,20,20,,,,,,
28,攻撃速度ⅡLv1,器用系統,パッシブ,攻撃速度を3%増加,4,12,,,,,,,,,,,,,,,,,,,
28,攻撃速度ⅡLv2,器用系統,パッシブ,攻撃速度を6%増加,5,36,10,,,,,,,,,,20,,,,,,,,
28,攻撃速度ⅡLv3,器用系統,パッシブ,攻撃速度を10%増加,6,96,20,,,,,,,,,,40,,,,,,,,
28,攻撃速度ⅡLv4,器用系統,パッシブ,攻撃速度を15%増加,7,168,40,,,,,,,,,,40,20,,,,,,,
28,攻撃速度ⅡLv5,器用系統,パッシブ,攻撃速度を20%増加,8,300,60,,,,,,,,,,40,20,20,,,,,,
317,魔法クリティカル発動率ⅠLv1,器用系統,パッシブ,魔法クリティカル発動率を3%増加,6,30,,,,,,,,,,,,,,,,,,,
317,魔法クリティカル発動率ⅠLv2,器用系統,パッシブ,魔法クリティカル発動率を6%増加,7,80,20,,,,,,,,,,40,,,,,,,,
317,魔法クリティカル発動率ⅠLv3,器用系統,パッシブ,魔法クリティカル発動率を10%増加,8,140,40,,,,,,,,,,40,20,,,,,,,
317,魔法クリティカル発動率ⅠLv4,器用系統,パッシブ,魔法クリティカル発動率を15%増加,9,250,80,,,,,,,,,,40,20,20,,,,,,
317,魔法クリティカル発動率ⅠLv5,器用系統,パッシブ,魔法クリティカル発動率を20%増加,10,400,120,,,,,,,,,,80,40,20,,,,,,
314,器用ⅡLv1,器用系統,パッシブ,器用を2%増加,7,30,,,,,,,,,,,,,,,,,,,
314,器用ⅡLv2,器用系統,パッシブ,器用を4%増加,8,80,20,,,,,,,,,,40,,,,,,,,
314,器用ⅡLv3,器用系統,パッシブ,器用を6%増加,9,140,40,,,,,,,,,,40,20,,,,,,,
314,器用ⅡLv4,器用系統,パッシブ,器用を10%増加,10,250,80,,,,,,,,,,40,20,20,,,,,,
314,器用ⅡLv5,器用系統,パッシブ,器用を15%増加,11,400,120,,,,,,,,,,80,40,20,,,,,,
316,物理クリティカル倍率Lv1,器用系統,パッシブ,物理クリティカル倍率を3%増加,8,30,,,,,,,,,,,,,,,,,,,
316,物理クリティカル倍率Lv2,器用系統,パッシブ,物理クリティカル倍率を6%増加,9,80,20,,,,,,,,,,40,,,,,,,,
316,物理クリティカル倍率Lv3,器用系統,パッシブ,物理クリティカル倍率を10%増加,10,140,40,,,,,,,,,,40,20,,,,,,,
316,物理クリティカル倍率Lv4,器用系統,パッシブ,物理クリティカル倍率を15%増加,11,250,80,,,,,,,,,,40,20,20,,,,,,
316,物理クリティカル倍率Lv5,器用系統,パッシブ,物理クリティカル倍率を20%増加,12,400,120,,,,,,,,,,80,40,20,,,,,,
315,専心Lv1,器用系統,アクティブ,180秒間、10秒毎にMPが1%ずつ回復。,10,50,50,,,,,,,,,,,,,,,,,,
315,専心Lv2,器用系統,アクティブ,180秒間、10秒毎にMPが2%ずつ回復。,11,100,100,,,,,,,,,,50,,,,,,,,
315,専心Lv3,器用系統,アクティブ,180秒間、10秒毎にMPが3%ずつ回復。,12,180,150,,,,,,,,,,60,30,,,,,,,
315,専心Lv4,器用系統,アクティブ,180秒間、10秒毎にMPが4%ずつ回復。,13,300,200,,,,,,,,,,70,40,20,,,,,,
315,専心Lv5,器用系統,アクティブ,180秒間、10秒毎にMPが5%ずつ回復。,14,450,250,,,,,,,,,,80,50,30,,,,,,
211,MPⅠLv1,精神系統,パッシブ,最大MPを2%増加,3,12,,,,,,,,,,,,,,,,,,,
211,MPⅠLv2,精神系統,パッシブ,最大MPを4%増加,4,36,10,,,,,,,,,,,,,,,,20,,
211,MPⅠLv3,精神系統,パッシブ,最大MPを6%増加,5,96,20,,,,,,,,,,,,,,,,40,,
211,MPⅠLv4,精神系統,パッシブ,最大MPを9%増加,6,168,40,,,,,,,,,,,,,,,,40,20,
211,MPⅠLv5,精神系統,パッシブ,最大MPを12%増加,7,300,60,,,,,,,,,,,,,,,,40,20,20
210,詠唱速度ⅠLv1,精神系統,パッシブ,詠唱速度を1.03倍する,4,12,,,,,,,,,,,,,,,,,,,
210,詠唱速度ⅠLv2,精神系統,パッシブ,詠唱速度を1.06倍する,5,36,10,,,,,,,,,,,,,,,,20,,
210,詠唱速度ⅠLv3,精神系統,パッシブ,詠唱速度を1.09倍する,6,96,20,,,,,,,,,,,,,,,,40,,
210,詠唱速度ⅠLv4,精神系統,パッシブ,詠唱速度を1.12倍する,7,168,40,,,,,,,,,,,,,,,,40,20,
210,詠唱速度ⅠLv5,精神系統,パッシブ,詠唱速度を1.15倍する,8,300,60,,,,,,,,,,,,,,,,40,20,20
321,魔法クリティカル発動率ⅡLv1,精神系統,パッシブ,魔法クリティカル発動率を3%増加,6,30,,,,,,,,,,,,,,,,,,,
321,魔法クリティカル発動率ⅡLv2,精神系統,パッシブ,魔法クリティカル発動率を6%増加,7,80,20,,,,,,,,,,,,,,,,40,,
321,魔法クリティカル発動率ⅡLv3,精神系統,パッシブ,魔法クリティカル発動率を10%増加,8,140,40,,,,,,,,,,,,,,,,40,20,
321,魔法クリティカル発動率ⅡLv4,精神系統,パッシブ,魔法クリティカル発動率を15%増加,9,250,80,,,,,,,,,,,,,,,,40,20,20
321,魔法クリティカル発動率ⅡLv5,精神系統,パッシブ,魔法クリティカル発動率を20%増加,10,400,120,,,,,,,,,,,,,,,,80,40,20
318,精神ⅡLv1,精神系統,パッシブ,精神を2%増加,8,30,,,,,,,,,,,,,,,,,,,
318,精神ⅡLv2,精神系統,パッシブ,精神を4%増加,9,80,20,,,,,,,,,,,,,,,,40,,
318,精神ⅡLv3,精神系統,パッシブ,精神を6%増加,10,140,40,,,,,,,,,,,,,,,,40,20,
318,精神ⅡLv4,精神系統,パッシブ,精神を10%増加,11,250,80,,,,,,,,,,,,,,,,40,20,20
318,精神ⅡLv5,精神系統,パッシブ,精神を15%増加,12,400,120,,,,,,,,,,,,,,,,80,40,20
320,魔法クリティカル倍率Lv1,精神系統,パッシブ,魔法クリティカル倍率を5%増加,7,30,,,,,,,,,,,,,,,,,,,
320,魔法クリティカル倍率Lv2,精神系統,パッシブ,魔法クリティカル倍率を7%増加,8,80,20,,,,,,,,,,,,,,,,40,,
320,魔法クリティカル倍率Lv3,精神系統,パッシブ,魔法クリティカル倍率を10%増加,9,140,40,,,,,,,,,,,,,,,,40,20,
320,魔法クリティカル倍率Lv4,精神系統,パッシブ,魔法クリティカル倍率を20%増加,10,250,80,,,,,,,,,,,,,,,,40,20,20
320,魔法クリティカル倍率Lv5,精神系統,パッシブ,魔法クリティカル倍率を30%増加,11,400,120,,,,,,,,,,,,,,,,80,40,20
319,求道Lv1,精神系統,アクティブ,HPが50%以下の時、魔法スキルの威力が10%アップする,10,50,50,,,,,,,,,,,,,,,,,,
319,求道Lv2,精神系統,アクティブ,HPが50%以下の時、魔法スキルの威力が20%アップする,11,100,100,,,,,,,,,,,,,,,,50,,
319,求道Lv3,精神系統,アクティブ,HPが50%以下の時、魔法スキルの威力が30%アップする,12,180,150,,,,,,,,,,,,,,,,60,30,
319,求道Lv4,精神系統,アクティブ,HPが50%以下の時、魔法スキルの威力が40%アップする,13,300,200,,,,,,,,,,,,,,,,70,40,20
319,求道Lv5,精神系統,アクティブ,HPが50%以下の時、魔法スキルの威力が50%アップする,14,450,250,,,,,,,,,,,,,,,,80,50,30